// lab61soc.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module lab61soc (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

endmodule
